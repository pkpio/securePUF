`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
// Author 			:	Praveen Kumar Pendyala
// Create Date		:  07/13/14
// Modify Date		:	07/13/14
// Module Name		:  pufInputNetwork
// Project Name   :  PDL
// Target Devices	: 	Xilinx Vertix 5, XUPV5 110T
// Tool versions	: 	14.4 ISE
//
// Description:
// This module does the XORing of challenges to satisfy the Strict Avalanche
//	Criterion (SAC) for a parallel PUF circuit as described in Lightweight Secure 
// PUFs paper.
//
//////////////////////////////////////////////////////////////////////////////////
module pufInputNetwork(
		
    );


endmodule
